module RX_element_VC0();


endmodule