module top();

endmodule